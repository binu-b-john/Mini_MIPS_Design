----------------------------------------------------------------------------------
-- Company: 	Concordia University
-- Engineer: 	Binu Basil John
-- 
-- Create Date:    21:23:26 09/10/2018 
-- Design Name: 
-- Module Name:    mini_MIPS - Behavioral 
-- Project Name:	 Mini_MIPS_Design
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity mini_MIPS is
    Port ( clk,rst : in  STD_LOGIC);
end mini_MIPS;

architecture Behavioral of mini_MIPS is

begin


end Behavioral;

